.option method=GEAR
.option accurate=1
*.option absv=1e-9 vfloor=1e-9 numdgt=10 ingold=1 lvltim=3 dvdt=3

* Standard.bjt models :

.MODEL BD139 NPN ( IS=2.3985E-13 BF=244.9 NF=1.0 BR=78.11 NR=1.007 ISE=1.0471E-14 NE=1.2 ISC=1.9314E-11 NC=1.45 VAF=98.5 VAR=7.46 IKF=1.1863 IKR=0.1445 RB=2.14 RBM=0.001 IRB=0.031 RE=0.0832 RC=0.01 CJE=2.92702E-10 VJE=0.67412 MJE=0.3300 FC=0.5 CJC=4.8831E-11 VJC=0.5258 MJC=0.3928 XCJC=0.5287 XTB=1.1398 EG=1.2105 XTI=3.0 Vceo=80 Icrating=3 mfg=fairchild )
.MODEL BD140 PNP ( IS=2.9537E-13 BF=201.4 NF=1.0 BR=23.765 NR=1.021 ISE=1.8002E-13 NE=1.5 ISC=7.0433p NC=1.38 VAF=137.0 VAR=8.41 IKF=1.0993 IKR=0.10 RB=1.98 RBM=0.01 IRB=0.011 RE=0.1109 RC=0.01 CJE=2.1982E-10 VJE=0.7211 MJE=0.3685 FC=0.5 CJC=6.8291E-11 VJC=0.5499 MJC=0.3668 XCJC=0.5287 XTB=1.4883 EG=1.2343 XTI=3.0 Vceo=80 Icrating=3 mfg=fairchild )
.MODEL BD135P NPN ( IS=4.815E-14 ISE=1.389E-14 ISC=1.295E-13 XTI=3 BF=124.2 BR=13.26 IKF=1.6 IKR=0.29 XTB=1.5 VAF=222 VAR=81.4 VJE=0.7313 VJC=0.5642 RE=0.165 RC=0.096 RB=0.5 RBM=0.5 IRB=1E-06 CJE=1.243E-10 CJC=3.04E-11 XCJC=0.15 FC=0.9359 NF=0.9897 NR=0.9895 NE=1.6 NC=1.183 MJE=0.3476 MJC=0.4371 TF=6.478E-10 TR=1m2 ITF=3.35 VTF=2.648 XTF=29 EG=1.11 VCEO=45 ICRATING=1.5 MFG=PHILIPS )
.MODEL BD136P PNP ( IS=7.401E-14 ISE=4.104E-16 ISC=1.290E-14 XTI=3 BF=336.5 BR=13.91 IKF=0.1689 IKR=9.888E-2 XTB=1.5 VAF=224.7 VAR=30.00 VJE=0.6900 VJC=0.6431 RE=0.208 RC=5.526E-02 RB=0.500 RBM=0.500 IRB=1E-06 CJE=1.066E-10 CJC=5.234E-11 XCJC=0.440 FC=0.990 NF=0.9938 NR=0.9913 NE=1.054 NC=1.100 MJE=0.3676 MJC=0.4436 TF=2.578E-10 TR=1E-25 ITF=1.3040 VTF=2.366 XTF=13.56 EG=1.11 VCEO=45 ICRATING=1.5 MFG=PHILIPS )

.model Q2N3904 NPN(IS=1E-14 VAF=100 Bf=300 IKF=0.4 XTB=1.5 BR=4 CJC=4E-12 CJE=8E-12 RB=20 RC=0.1 RE=0.1 TR=250E-9 TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)
.model Q2N3906 PNP(IS=1E-14 VAF=100 BF=200 IKF=0.4 XTB=1.5 BR=4 CJC=4.5E-12 CJE=10E-12 RB=20 RC=0.1 RE=0.1 TR=250E-9 TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)

.model D1N4148  D 
+Is=2.682n N=1.836 Rs=.5664 Xti=3 Eg=1.11 Cjo=4p
+M=.3333 Vj=.5 Fc=.5 Bv=100 Ibv=100u Tt=11.54n

.model Dbreak D Is=1e-14 Cjo=.1pF Rs=.1 BV=5V IBV=2mA

*********************************Netlist**************************
* Sources
VCC     	200		0  		15
VEE		100		0		-15
*VIN1		1		0		sin(0	141.4m	1k	0	0)
VIN		1		0		AC		1

** Buffer Stage
R1		2		100		15.6693k
Rx1		200		2		14.3307k
Rx2		3		100		15k		

Qx1		200		2		3		Q2N3904

C4		1		2		2.2u

** Differential Ampilifier
R2		5		100		7.15k
R3		4		12		1x
RBQ2		4		0		10

C1		4		0		100p
C2		22		0		47u

Q1		6		3		5		Q2N3904
Q2		7		4		5		Q2N3904
Q8		10		8		7		Q2N3904
Q9		9		8		6		Q2N3904
Q6		10		9		200		Q2N3906
Q7		9		9		200		Q2N3906

Vb		8		0		2

** Z
Qz		13		11		12		Q2N3904

Rz1		200		11		13k
Rz2		11		0		2k

Rz3		12		0		1k
Rz4		200		13		5k

C3		13		15		100p
R		10		11		0

*Cz		10		11		100u
*Dz		10		0		Dbreak
*Rbias1		10		500		1k
*Rbias2		10		100		200

** Output Stage
R4		17		100		3k
R6		18		19		1
R7		19		20		1
RL		21		0		8
RCQ3		14		200		1.45k

Q3		15		13		14		Q2N3906
Q4		200		15		18		Q2N3904
Q5		100		17		20		Q2N3906

CL		19		21		100m

D1		15		16		D1N4148
D2		16		17		D1N4148

** FeedBack
RF		21		4		143

******************************************************************
.op
*.TRAN	1us	10ms
*.AC DEC 40 1 20k
.AC LIN 100 1 100
.end

